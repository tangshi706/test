module test(input clk,input rst_n,input a,input b,input cin,output sum,output co);

assign {co,sum}=a+b+ci;

endmodule 
